module module1();
endmodule
